all rtl design file
