all testbench component files
